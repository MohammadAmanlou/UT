`timescale 1ns/1ns
module Q1Nand(input a , b , output w);
	supply1 Vdd;
	supply0 Gnd;
	wire y;
	pmos #(5,6,7) P1(w,Vdd,a) , P2(w,Vdd,b);
	nmos #(3,4,5) N1(y,Gnd,b) , N2(w,y,a);
endmodule