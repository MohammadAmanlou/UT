`timescale 1ns/1ns
module ALU_2(input [7:0]a,b,input[2:0]f,output [7:0]w,output c,output z);
	wire s;
	reg cin=1'b0;
	reg [7:0]bsel,m;
	wire [7:0] sum;
	CRA_8bit adder(a,bsel,cin,sum,c);
	assign bsel=(f[1]&f[0])?b>>1:
  		(~f[1]&f[0])?b<<1:
  		(~f[1]&~f[0])?b:8'b0;
	assign s=sum[7];
	assign m=(f[1]&~f[0]&s)?b:
   		(f[1]&~f[0]&~s)?a:
  		(~(f[1]&~f[0]))?sum:8'b0;
	assign en=f[2]&~f[1]&~f[0];
	assign w=en?8'b0:
  		(f[2]==1'b0)?m:
  		(f==3'b100)?8'b0:
  		(f==3'b101)?a|b:
  		(f==3'b110)?a&b:
  		(f==3'b111)?b<<1:8'b0;
	assign z=~|w;
endmodule
