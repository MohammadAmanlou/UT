module Adder(
  input [8:0] A,
  input [8:0] B,
  output [8:0] Sum
);


  assign Sum = A + B ;


endmodule
